module Mealy(
 din,
 clk,
reset,
 y
    );
input din,clk,reset;
output reg y;
parameter S0=3'b000, S1=3'b001, S2=3'b010, S3=3'b011, S4=3'b100, S5=3'b101;
reg [2:0]nextState;
always @(posedge clk)
begin
if(reset)
begin
y=0;
nextState=S0;
end
else
case(nextState)
S0:
begin
if(din==0)
begin
nextState=S1;
y=0;
end
else
begin
nextState=S0;
y=0;
end
end
S1:
begin
if(din==0)
begin
nextState=S3;
y=0;
end
else
begin
nextState=S2;
y=0;
end
end
S2:
begin
if(din==0)
begin
nextState=S5;
y=0;
end
else
begin
nextState=S0;
y=0;
end
end
S3:
begin
if(din==0)
begin
nextState=S4;
y=0;
end
else
begin
nextState=S2;
y=0;
end
end
S4:
begin
if(din==0)
begin
nextState=S4;
y=0;
end
else
begin
nextState=S2;
y=1;
end
end
S5:
begin
if(din==0)
begin
nextState=S3;
y=0;
end
else
begin
nextState=S2;
y=1;
end
end
endcase
end
endmodule
